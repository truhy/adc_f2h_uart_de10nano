// soc_system.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                         //                 clk.clk
		input  wire        hps_0_f2h_axi_clock_clk,         // hps_0_f2h_axi_clock.clk
		input  wire [7:0]  hps_0_f2h_axi_slave_awid,        // hps_0_f2h_axi_slave.awid
		input  wire [31:0] hps_0_f2h_axi_slave_awaddr,      //                    .awaddr
		input  wire [3:0]  hps_0_f2h_axi_slave_awlen,       //                    .awlen
		input  wire [2:0]  hps_0_f2h_axi_slave_awsize,      //                    .awsize
		input  wire [1:0]  hps_0_f2h_axi_slave_awburst,     //                    .awburst
		input  wire [1:0]  hps_0_f2h_axi_slave_awlock,      //                    .awlock
		input  wire [3:0]  hps_0_f2h_axi_slave_awcache,     //                    .awcache
		input  wire [2:0]  hps_0_f2h_axi_slave_awprot,      //                    .awprot
		input  wire        hps_0_f2h_axi_slave_awvalid,     //                    .awvalid
		output wire        hps_0_f2h_axi_slave_awready,     //                    .awready
		input  wire [4:0]  hps_0_f2h_axi_slave_awuser,      //                    .awuser
		input  wire [7:0]  hps_0_f2h_axi_slave_wid,         //                    .wid
		input  wire [31:0] hps_0_f2h_axi_slave_wdata,       //                    .wdata
		input  wire [3:0]  hps_0_f2h_axi_slave_wstrb,       //                    .wstrb
		input  wire        hps_0_f2h_axi_slave_wlast,       //                    .wlast
		input  wire        hps_0_f2h_axi_slave_wvalid,      //                    .wvalid
		output wire        hps_0_f2h_axi_slave_wready,      //                    .wready
		output wire [7:0]  hps_0_f2h_axi_slave_bid,         //                    .bid
		output wire [1:0]  hps_0_f2h_axi_slave_bresp,       //                    .bresp
		output wire        hps_0_f2h_axi_slave_bvalid,      //                    .bvalid
		input  wire        hps_0_f2h_axi_slave_bready,      //                    .bready
		input  wire [7:0]  hps_0_f2h_axi_slave_arid,        //                    .arid
		input  wire [31:0] hps_0_f2h_axi_slave_araddr,      //                    .araddr
		input  wire [3:0]  hps_0_f2h_axi_slave_arlen,       //                    .arlen
		input  wire [2:0]  hps_0_f2h_axi_slave_arsize,      //                    .arsize
		input  wire [1:0]  hps_0_f2h_axi_slave_arburst,     //                    .arburst
		input  wire [1:0]  hps_0_f2h_axi_slave_arlock,      //                    .arlock
		input  wire [3:0]  hps_0_f2h_axi_slave_arcache,     //                    .arcache
		input  wire [2:0]  hps_0_f2h_axi_slave_arprot,      //                    .arprot
		input  wire        hps_0_f2h_axi_slave_arvalid,     //                    .arvalid
		output wire        hps_0_f2h_axi_slave_arready,     //                    .arready
		input  wire [4:0]  hps_0_f2h_axi_slave_aruser,      //                    .aruser
		output wire [7:0]  hps_0_f2h_axi_slave_rid,         //                    .rid
		output wire [31:0] hps_0_f2h_axi_slave_rdata,       //                    .rdata
		output wire [1:0]  hps_0_f2h_axi_slave_rresp,       //                    .rresp
		output wire        hps_0_f2h_axi_slave_rlast,       //                    .rlast
		output wire        hps_0_f2h_axi_slave_rvalid,      //                    .rvalid
		input  wire        hps_0_f2h_axi_slave_rready,      //                    .rready
		output wire        hps_0_h2f_reset_reset_n,         //     hps_0_h2f_reset.reset_n
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //              hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //                    .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //                    .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //                    .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //                    .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //                    .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //                    .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //                    .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //                    .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //                    .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //                    .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //                    .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //                    .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //                    .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //                    .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //                    .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //                    .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //                    .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //                    .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //                    .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //                    .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //                    .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //                    .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //                    .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //                    .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //                    .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //                    .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //                    .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //                    .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //                    .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //                    .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //                    .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,    //                    .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,   //                    .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,   //                    .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,    //                    .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,     //                    .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //                    .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,     //                    .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,     //                    .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,     //                    .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,     //                    .hps_io_i2c1_inst_SCL
		output wire [14:0] memory_mem_a,                    //              memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //                    .mem_ba
		output wire        memory_mem_ck,                   //                    .mem_ck
		output wire        memory_mem_ck_n,                 //                    .mem_ck_n
		output wire        memory_mem_cke,                  //                    .mem_cke
		output wire        memory_mem_cs_n,                 //                    .mem_cs_n
		output wire        memory_mem_ras_n,                //                    .mem_ras_n
		output wire        memory_mem_cas_n,                //                    .mem_cas_n
		output wire        memory_mem_we_n,                 //                    .mem_we_n
		output wire        memory_mem_reset_n,              //                    .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //                    .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //                    .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //                    .mem_dqs_n
		output wire        memory_mem_odt,                  //                    .mem_odt
		output wire [3:0]  memory_mem_dm,                   //                    .mem_dm
		input  wire        memory_oct_rzqin,                //                    .oct_rzqin
		output wire        pll_0_locked_export,             //        pll_0_locked.export
		output wire        pll_0_outclk0_clk,               //       pll_0_outclk0.clk
		output wire        pll_0_outclk1_clk,               //       pll_0_outclk1.clk
		input  wire        reset_reset_n                    //               reset.reset_n
	);

	soc_system_hps_0 #(
		.F2S_Width (1),
		.S2F_Width (0)
	) hps_0 (
		.mem_a                    (memory_mem_a),                    //        memory.mem_a
		.mem_ba                   (memory_mem_ba),                   //              .mem_ba
		.mem_ck                   (memory_mem_ck),                   //              .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                 //              .mem_ck_n
		.mem_cke                  (memory_mem_cke),                  //              .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                 //              .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                //              .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                //              .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                 //              .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),              //              .mem_reset_n
		.mem_dq                   (memory_mem_dq),                   //              .mem_dq
		.mem_dqs                  (memory_mem_dqs),                  //              .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                //              .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                  //              .mem_odt
		.mem_dm                   (memory_mem_dm),                   //              .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                //              .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK), //        hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),   //              .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),   //              .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),   //              .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),   //              .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),   //              .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),   //              .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),    //              .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL), //              .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL), //              .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK), //              .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),   //              .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),   //              .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),   //              .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),     //              .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),      //              .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),      //              .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),     //              .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),      //              .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),      //              .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),      //              .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),      //              .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),      //              .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),      //              .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),      //              .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),      //              .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),      //              .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),      //              .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),     //              .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),     //              .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),     //              .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),     //              .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),    //              .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),   //              .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),   //              .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),    //              .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),     //              .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),     //              .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),     //              .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),     //              .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),     //              .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),     //              .hps_io_i2c1_inst_SCL
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),         //     h2f_reset.reset_n
		.f2h_axi_clk              (hps_0_f2h_axi_clock_clk),         // f2h_axi_clock.clk
		.f2h_AWID                 (hps_0_f2h_axi_slave_awid),        // f2h_axi_slave.awid
		.f2h_AWADDR               (hps_0_f2h_axi_slave_awaddr),      //              .awaddr
		.f2h_AWLEN                (hps_0_f2h_axi_slave_awlen),       //              .awlen
		.f2h_AWSIZE               (hps_0_f2h_axi_slave_awsize),      //              .awsize
		.f2h_AWBURST              (hps_0_f2h_axi_slave_awburst),     //              .awburst
		.f2h_AWLOCK               (hps_0_f2h_axi_slave_awlock),      //              .awlock
		.f2h_AWCACHE              (hps_0_f2h_axi_slave_awcache),     //              .awcache
		.f2h_AWPROT               (hps_0_f2h_axi_slave_awprot),      //              .awprot
		.f2h_AWVALID              (hps_0_f2h_axi_slave_awvalid),     //              .awvalid
		.f2h_AWREADY              (hps_0_f2h_axi_slave_awready),     //              .awready
		.f2h_AWUSER               (hps_0_f2h_axi_slave_awuser),      //              .awuser
		.f2h_WID                  (hps_0_f2h_axi_slave_wid),         //              .wid
		.f2h_WDATA                (hps_0_f2h_axi_slave_wdata),       //              .wdata
		.f2h_WSTRB                (hps_0_f2h_axi_slave_wstrb),       //              .wstrb
		.f2h_WLAST                (hps_0_f2h_axi_slave_wlast),       //              .wlast
		.f2h_WVALID               (hps_0_f2h_axi_slave_wvalid),      //              .wvalid
		.f2h_WREADY               (hps_0_f2h_axi_slave_wready),      //              .wready
		.f2h_BID                  (hps_0_f2h_axi_slave_bid),         //              .bid
		.f2h_BRESP                (hps_0_f2h_axi_slave_bresp),       //              .bresp
		.f2h_BVALID               (hps_0_f2h_axi_slave_bvalid),      //              .bvalid
		.f2h_BREADY               (hps_0_f2h_axi_slave_bready),      //              .bready
		.f2h_ARID                 (hps_0_f2h_axi_slave_arid),        //              .arid
		.f2h_ARADDR               (hps_0_f2h_axi_slave_araddr),      //              .araddr
		.f2h_ARLEN                (hps_0_f2h_axi_slave_arlen),       //              .arlen
		.f2h_ARSIZE               (hps_0_f2h_axi_slave_arsize),      //              .arsize
		.f2h_ARBURST              (hps_0_f2h_axi_slave_arburst),     //              .arburst
		.f2h_ARLOCK               (hps_0_f2h_axi_slave_arlock),      //              .arlock
		.f2h_ARCACHE              (hps_0_f2h_axi_slave_arcache),     //              .arcache
		.f2h_ARPROT               (hps_0_f2h_axi_slave_arprot),      //              .arprot
		.f2h_ARVALID              (hps_0_f2h_axi_slave_arvalid),     //              .arvalid
		.f2h_ARREADY              (hps_0_f2h_axi_slave_arready),     //              .arready
		.f2h_ARUSER               (hps_0_f2h_axi_slave_aruser),      //              .aruser
		.f2h_RID                  (hps_0_f2h_axi_slave_rid),         //              .rid
		.f2h_RDATA                (hps_0_f2h_axi_slave_rdata),       //              .rdata
		.f2h_RRESP                (hps_0_f2h_axi_slave_rresp),       //              .rresp
		.f2h_RLAST                (hps_0_f2h_axi_slave_rlast),       //              .rlast
		.f2h_RVALID               (hps_0_f2h_axi_slave_rvalid),      //              .rvalid
		.f2h_RREADY               (hps_0_f2h_axi_slave_rready)       //              .rready
	);

	soc_system_pll_0 pll_0 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),   // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk),   // outclk1.clk
		.locked   (pll_0_locked_export)  //  locked.export
	);

endmodule
